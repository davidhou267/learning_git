module test_git (
    input   clk,
    input   rst_n,
    input   data_in,
    output  data_out
);
    
endmodule