module test_git (
    input   clk,
    input   rst_n
);
    
endmodule